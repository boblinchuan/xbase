{{ _header }}

// Intentionally nothing, since this does nothing logically.

endmodule
